`define FPGA

//`define OPENLANE

`ifdef OPENLANE
    `define GATE _sky130
`else
    `define GATE
`endif


// Parameters
`define DATA_WIDTH 32
`define REG_DATA_WIDTH 32   // Word Width
`define REG_ADDR_WIDTH 5   // Address With
`define REG_DEPTH 1 << `REG_ADDR_WIDTH  // Total number of positions (32)


`define MEM_DATA_WIDTH 32   // Word Width
`define MEM_ADDR_WIDTH 10   // Address With
`define MEM_DEPTH 1 << `MEM_ADDR_WIDTH-2  // Total number of positions (1024)

`define MEM_TRANSFER_WIDTH 4  // Mask to store word, halfword or byte


// RV32IM Buyruklari

`define ADD        32'b0000000??????????000?????0110011
`define ADDI       32'b?????????????????000?????0010011
`define AND        32'b0000000??????????111?????0110011
`define ANDI       32'b?????????????????111?????0010011
`define AUIPC      32'b?????????????????????????0010111
`define BEQ        32'b?????????????????000?????1100011
`define BGE        32'b?????????????????101?????1100011
`define BGEU       32'b?????????????????111?????1100011
`define BLT        32'b?????????????????100?????1100011
`define BLTU       32'b?????????????????110?????1100011
`define BNE        32'b?????????????????001?????1100011
`define DIV        32'b0000001??????????100?????0110011
`define DIVU       32'b0000001??????????101?????0110011
`define EBREAK     32'b00000000000100000000000001110011
`define ECALL      32'b00000000000000000000000001110011
`define FENCE      32'b?????????????????000?????0001111
`define FENCE_I    32'b?????????????????001?????0001111
`define JAL        32'b?????????????????????????1101111
`define JALR       32'b?????????????????000?????1100111
`define LB         32'b?????????????????000?????0000011
`define LBU        32'b?????????????????100?????0000011
`define LH         32'b?????????????????001?????0000011
`define LHU        32'b?????????????????101?????0000011
`define LUI        32'b?????????????????????????0110111
`define LW         32'b?????????????????010?????0000011
`define MUL        32'b0000001??????????000?????0110011
`define MULH       32'b0000001??????????001?????0110011
`define MULHSU     32'b0000001??????????010?????0110011
`define MULHU      32'b0000001??????????011?????0110011
`define OR         32'b0000000??????????110?????0110011
`define ORI        32'b?????????????????110?????0010011
`define REM        32'b0000001??????????110?????0110011
`define REMU       32'b0000001??????????111?????0110011
`define SB         32'b?????????????????000?????0100011
`define SH         32'b?????????????????001?????0100011
`define SLL        32'b0000000??????????001?????0110011
`define SLLI       32'b0000000??????????001?????0010011
`define SLT        32'b0000000??????????010?????0110011
`define SLTI       32'b?????????????????010?????0010011
`define SLTIU      32'b?????????????????011?????0010011
`define SLTU       32'b0000000??????????011?????0110011
`define SRA        32'b0100000??????????101?????0110011
`define SRAI       32'b0100000??????????101?????0010011
`define SRL        32'b0000000??????????101?????0110011
`define SRLI       32'b0000000??????????101?????0010011
`define SUB        32'b0100000??????????000?????0110011
`define SW         32'b?????????????????010?????0100011
`define XOR        32'b0000000??????????100?????0110011
`define XORI       32'b?????????????????100?????0010011



// RV32A Buyruklari

`define LR_W        32'b00010??????????010?????0101111
`define SC_W        32'b00011??????????010?????0101111
`define AMOSWAP_W   32'b00001??????????010?????0101111
`define AMOADD_W    32'b00000??????????010?????0101111
`define AMOXOR_W    32'b00100??????????010?????0101111
`define AMOAND_W    32'b01100??????????010?????0101111
`define AMOOR_W     32'b01000??????????010?????0101111
`define AMOMIN_W    32'b10000??????????010?????0101111
`define AMOMAX_W    32'b10100??????????010?????0101111
`define AMOMINU_W   32'b11000??????????010?????0101111
`define AMOMAXU_W   32'b11100??????????010?????0101111

/*
// RV32F Buyruklari
`define FLW         32'b?????????????????010?????0000111
`define FSW         32'b?????????????????010?????0100111
`define FMADD_S     32'b?????00??????????000?????1000011
`define FMSUB_S     32'b?????00??????????000?????1000111
`define FNMSUB_S    32'b?????00??????????000?????1001011
`define FNMADD_S    32'b?????00??????????000?????1001111
`define FADD_S      32'b0000000??????????000?????1010011
`define FSUB_S      32'b0000100??????????000?????1010011
`define FMUL_S      32'b0001000??????????000?????1010011
`define FDIV_S      32'b0001100??????????000?????1010011
`define FSQRT_S     32'b010110000000?????000?????1010011
`define FSGNJ_S     32'b0010000??????????000?????1010011
`define FSGNJN_S    32'b0010000??????????001?????1010011
`define FSGNJX_S    32'b0010000??????????010?????1010011
`define FMIN_S      32'b0010100??????????000?????1010011
`define FMAX_S      32'b0010100??????????001?????1010011
`define FCVT_W_S    32'b110000000000?????000?????1010011
`define FCVT_WU_S   32'b110000000001?????000?????1010011
`define FMV_X_W     32'b111000000000?????000?????1010011
`define FEQ_S       32'b1010000??????????010?????1010011
`define FLT_S       32'b1010000??????????001?????1010011
`define FLE_S       32'b1010000??????????000?????1010011
`define FCLASS_S    32'b111000000000?????001?????1010011
`define FCVT_S_W    32'b110100000000?????000?????1010011 
`define FCVT_S_WU   32'b110100000001?????000?????1010011
`define FMV_W_X     32'b111100000000?????000?????1010011
*/

// RV32B Buyruklari

// rvb_zbb32_macros.vh

`define INSN_OPNEG_ANDN  32'b0100000??????????111?????0110011
`define INSN_OPNEG_ORN   32'b0100000??????????110?????0110011
`define INSN_OPNEG_XNOR  32'b0100000??????????100?????0110011
`define INSN_SHIFT_SLL   32'b0000000??????????001?????0110011
`define INSN_SHIFT_SRL   32'b0000000??????????101?????0110011
`define INSN_SHIFT_SRA   32'b0100000??????????101?????0110011
`define INSN_SHIFT_SLO   32'b0010000??????????001?????0110011
`define INSN_SHIFT_SRO   32'b0010000??????????101?????0110011
`define INSN_SHIFT_ROL   32'b0110000??????????001?????0110011
`define INSN_SHIFT_ROR   32'b0110000??????????101?????0110011
`define INSN_SHIFT_REV   32'b011010011111?????101?????0010011
`define INSN_SHIFT_REV8  32'b011010011000?????101?????0010011
`define INSN_SHIFT_ORC_B 32'b001010000111?????101?????0010011
`define INSN_BITCNT_CLZ  32'b011000000000?????001?????0010011
`define INSN_BITCNT_CTT  32'b011000000001?????001?????0010011
`define INSN_BITCNT_PCNT 32'b011000000010?????001?????0010011
`define INSN_MINMAX_MIN  32'b0000101??????????100?????0110011
`define INSN_MINMAX_MAX  32'b0000101??????????101?????0110011
`define INSN_MINMAX_MINU 32'b0000101??????????110?????0110011
`define INSN_MINMAX_MAXU 32'b0000101??????????111?????0110011
`define INSN_PACK        32'b0000100??????????100?????0110011

/*
`define ANDN        32'b0100000??????????111?????0110011
`define XNOR        32'b0100000??????????100?????0110011
`define SLO         32'b0010000??????????001?????0110011
`define SRO         32'b0010000??????????101?????0110011
`define ROL         32'b0110000??????????001?????0110011
`define ROR         32'b0110000??????????101?????0110011
`define SH1ADD      32'b0010000??????????010?????0110011
`define SH2ADD      32'b0010000??????????100?????0110011
`define SH3ADD      32'b0010000??????????110?????0110011
`define SBCLR       32'b0100100??????????001?????0110011
`define SBSET       32'b0010100??????????001?????0110011
`define SBINV       32'b0110100??????????001?????0110011
`define SBEXT       32'b0100100??????????101?????0110011
`define GORC        32'b0010100??????????101?????0110011
`define GREV        32'b0110100??????????101?????0110011
`define CMIX        32'b0000101??????????001?????0110011
`define CMOV        32'b0000101??????????101?????0110011
`define FSR         32'b0000100??????????101?????0110011 
`define CRC32_B     32'b1101000??????????100?????0110011
`define CRC32_H     32'b1101000??????????101?????0110011 
`define CRC32_W     32'b1101000??????????110?????0110011
`define CRC32C_B    32'b1101000??????????110?????0110011 
`define CRC32C_H    32'b1101100??????????101?????0110011
`define CRC32C_W    32'b1101100??????????110?????0110011 
`define CLMUL       32'b0000101??????????001?????0110011
`define CLMULR      32'b0000101??????????010?????0110011 
`define CLMULH      32'b0000101??????????011?????0110011
`define MIN         32'b0000101??????????100?????0110011 
`define MAX         32'b0000101??????????101?????0110011
`define MINU        32'b0000101??????????110?????0110011 
`define MAXU        32'b0000101??????????111?????0110011
`define BDEP        32'b0000100??????????110?????0110011 
`define BEXT        32'b0000100??????????111?????0110011
`define PACK        32'b0000100??????????100?????0110011 
`define PACKU       32'b0100100??????????100?????0110011
`define PACKH       32'b0000100??????????111?????0110011
`define CLZ         32'b0110000??????????001?????0010011 // Count Leading Zeros
`define CPOP        32'b0110000??????????001?????0010011 // Count Population (Set Bits)
`define CTZ         32'b0110000??????????001?????0010011 // Count Trailing Zeros
`define ORC         32'b0010100??????????101?????0010011 // Bitwise OR with Complement
`define ORN         32'b0100000??????????110?????0110011 // Bitwise OR with Inverted operand
`define REV8        32'b0110100??????????101?????0010011 // Byte-wise Reverse
`define RORI        32'b0110000??????????101?????0010011 // Rotate Right Immediate
`define BCLR        32'b0100100??????????001?????0110011 // Bit Clear
`define BCLRI       32'b0100100??????????001?????0010011 // Bit Clear Immediate
`define BEXTI       32'b0000100??????????110?????0010011 // Bit Extract Immediate
`define BINVI       32'b0110100??????????001?????0010011 // Bit Invert Immediate
`define BSETI       32'b0010100??????????001?????0010011 // Bit Set Immediate
`define SEXT_B      32'b0110000??????????000?????0010011 // Sign-extend Byte
`define SEXT_H      32'b0110000??????????001?????0010011 // Sign-extend Halfword
`define ZEXT_H      32'b0110000??????????010?????0010011 // Zero-extend Halfword
*/

// Buyruklarin cozulmesi icin gereken bitler 14 bit
// 30:29, 27, 25, 21:20, 14:12, 6:2
`define BUYRUK_COZ_BIT 14

`define EBREAK_COZ      14'b00000100011100
`define ECALL_COZ       14'b00000000011100
`define ADD_COZ         14'b0000??00001100
`define AND_COZ         14'b0000??11101100
`define DIV_COZ         14'b0001??10001100
`define DIVU_COZ        14'b0001??10101100
`define MUL_COZ         14'b0001??00001100
`define MULH_COZ        14'b0001??00101100
`define MULHSU_COZ      14'b0001??01001100
`define MULHU_COZ       14'b0001??01101100
`define OR_COZ          14'b0000??11001100
`define REM_COZ         14'b0001??11001100
`define REMU_COZ        14'b0001??11101100
`define SLL_COZ         14'b0000??00101100
`define SLT_COZ         14'b0000??01001100
`define SLTU_COZ        14'b0000??01101100
`define SRA_COZ         14'b1000??10101100
`define SRL_COZ         14'b0000??10101100
`define SUB_COZ         14'b1000??00001100
`define XOR_COZ         14'b0000??10001100
`define SLADD_COZ       14'b0100??01001100
`define SLLI_COZ        14'b000???00100100
`define SRAI_COZ        14'b100???10100100
`define SRLI_COZ        14'b000???10100100
`define ADDI_COZ        14'b??????00000100
`define ANDI_COZ        14'b??????11100100
`define BEQ_COZ         14'b??????00011000
`define BGE_COZ         14'b??????10111000
`define BGEU_COZ        14'b??????11111000
`define BLT_COZ         14'b??????10011000
`define BLTU_COZ        14'b??????11011000
`define BNE_COZ         14'b??????00111000
`define FENCE_COZ       14'b??????00000011
`define FENCE_I_COZ     14'b??????00100011
`define JALR_COZ        14'b??????00011001
`define LB_COZ          14'b??????00000000
`define LBU_COZ         14'b??????10000000
`define LH_COZ          14'b??????00100000
`define LHU_COZ         14'b??????10100000
`define LW_COZ          14'b??????01000000
`define ORI_COZ         14'b??????11000100
`define SB_COZ          14'b??????00001000
`define SH_COZ          14'b??????00101000
`define SLTI_COZ        14'b??????01000100
`define SLTIU_COZ       14'b??????01100100
`define SW_COZ          14'b??????01001000
`define XORI_COZ        14'b??????10000100
`define AUIPC_COZ       14'b?????????00101
`define JAL_COZ         14'b?????????11011
`define LUI_COZ         14'b?????????01101


`define LRW_COZ         14'b00010??0?01001
`define SCW_COZ         14'b00011????01001
`define AMOSWAP_COZ     14'b00001????01001
`define AMOADD_COZ      14'b00000????01001
`define AMOXOR_COZ      14'b00100????01001
`define AMOAND_COZ      14'b01100????01001
`define AMOOR_COZ       14'b10000????01001
`define AMOMIN_COZ      14'b00100????01001
`define AMOMAX_COZ      14'b10100????01001
`define AMOMINU_COZ     14'b11000????01001
`define AMOMAXU_COZ     14'b11100????01001



// Mikroislemler
`define MI_BIT 28

`define GERIYAZ   01:00
`define YAZMAC    02:02
`define OPERAND   04:03
`define BIRIM     07:05
`define DAL       10:08
`define ALU       14:11
`define BOLME     16:15
`define CARPMA    18:17
`define BIB       21:19


`define GERIYAZ_KAYNAK_YOK    2'd0
`define GERIYAZ_KAYNAK_YURUT  2'd1
`define GERIYAZ_KAYNAK_PC     2'd2
`define GERIYAZ_KAYNAK_CARP   2'd3

`define YAZMAC_YAZMA 1'b0
`define YAZMAC_YAZ   1'b1

`define OPERAND_REG      2'b00
`define OPERAND_IMM      2'b01
`define OPERAND_PC       2'b10
`define OPERAND_PCIMM    2'b11

`define BIRIM_ALU        3'h0
`define BIRIM_CARPMA     3'h1
`define BIRIM_BOLME      3'h2
`define BIRIM_BIB        3'h3
`define BIRIM_SISTEM     3'h4

`define DAL_EQ     3'b000
`define DAL_NE     3'b001
`define DAL_LT     3'b010
`define DAL_GE     3'b011
`define DAL_LTU    3'b100
`define DAL_GEU    3'b101
`define DAL_JAL    3'b110
`define DAL_JALR   3'b110
`define DAL_YOK    3'b111

//----Dallanma �ng�r�c� Tanimlamalar----
`define BTB_SATIR_SAYISI         32
`define BTB_PS_BIT               5
`define BTB_SATIR_BOYUT          (32 - `BTB_PS_BIT) + 1 + 32
`define BHT_SATIR_SAYISI         32
`define BHT_PS_BIT               5
`define DALLANMA_TAHMIN_BIT      2 // ilerde �ift kutuplu yap�labilir
`define BHT_SATIR_BOYUT          (32 - `BHT_PS_BIT) + `DALLANMA_TAHMIN_BIT
`define GENEL_GECMIS_YAZMACI_BIT 5
`define BTB_VALID_BITI           `BTB_SATIR_BOYUT-1 // en anlaml� biti
`define GGY_SAYAC_BIT            3



`define ALU_TOPLAMA  4'h0
`define ALU_CIKARMA  4'h1
`define ALU_XOR      4'h2
`define ALU_OR       4'h3
`define ALU_AND      4'h4
`define ALU_SLL      4'h5
`define ALU_SRL      4'h6
`define ALU_SRA      4'h7
`define ALU_SLT      4'h8
`define ALU_SLTU     4'h9
`define ALU_GECIR    4'ha
`define ALU_YOK      4'h0

`define BOLME_DIVU  2'h0
`define BOLME_REMU  2'h1
`define BOLME_DIV   2'h2
`define BOLME_REM   2'h3
`define BOLME_YOK   2'h0

`define CARPMA_MUL    2'h0
`define CARPMA_MULH   2'h1
`define CARPMA_MULHSU 2'h2
`define CARPMA_MULHU  2'h3
`define CARPMA_YOK    2'h0

// ALU_F OP-FP {funct7[6:2]};
`define FPU_FADD       5'b00000
`define FPU_FSUB       5'b00001
`define FPU_FMUL       5'b00010
`define FPU_FDIV       5'b00011
`define FPU_FSQRT      5'b01011
`define FPU_FSGNJ      5'b00100 // FSGNJ, FSGNJN, FSGNJX use rm to differentiate
`define FPU_FMINMAX    5'b00101 // FMIN, FMAX use rm to differentiate
`define FPU_FCVT_W_F   5'b11000 // FCVT.W/WU.S/L/D/Q
`define FPU_FMV_X      5'b11100 // also FCLASS, which uses rm to differentiate
`define FPU_FEQ        5'b10100 // FEQ, FLT, FLE use rm to differentiate
`define FPU_FCVT_F_W   5'b11010 // FCVT.S/L/D/Q.W and FCVT.S/L/D/Q.WU uses rm to diff
`define FPU_FMV_W_X    5'b11110

// FPU_F Fused Operations {2'b10, opcode[4:2]}
`define FPU_FMADD      5'b10000
`define FPU_FMSUB      5'b10001
`define FPU_FNMSUB     5'b10010
`define FPU_FNMADD     5'b10011

// FCSR
`define FRM_RNE 3'b000 // Round to Nearest, ties to Even
`define FRM_RTZ 3'b001 // Rounds towards Zero
`define FRM_RDN 3'b010 // Rounds Down (towards -inf)
`define FRM_RUP 3'b011 // Rounds Up (towards +inf)
`define FRM_RMM 3'b100 // Round to Nearest, ties to Max Magnitude
`define FRM_DYN 3'b111 // Use FCSR rounding mode

`define BIB_LB        3'h0
`define BIB_LBU       3'h1
`define BIB_LH        3'h2
`define BIB_LHU       3'h3
`define BIB_LW        3'h4
`define BIB_SB        3'h5
`define BIB_SH        3'h6
`define BIB_SW        3'h7
`define BIB_YOK       3'h0


// Diger SABITLER

// Buyruk tipleri
`define I_Tipi   3'b000
`define S_Tipi   3'b001
`define R_Tipi   3'b010
`define U_Tipi   3'b011
`define J_Tipi   3'b100
`define B_Tipi   3'b101
`define SYS_Tipi 3'b110

// DDB sabitleri
`define YON_GERIYAZ  2'b00
`define YON_YURUT    2'b01
`define YON_YOK      2'b10

// Dallanma Ongorucu Sabitleri
`define YANLIS_ATLADI 2'd3
`define ATLAMAMALIYDI 2'd2
`define ATLAMALIYDI   2'd1
`define SORUN_YOK     2'd0
// SORUN_YOK 0 olmak zorunda.

//-----------Bellek---------------
`define ADRES_BIT           32
`define BELLEK_BASLANGIC    32'h4000_0000
`define BELLEK_BOYUT        32'h0004_0000

//-----------Adres Aral�klar�-----------
`define UART_BASE_ADDR      32'h2000_0000
`define UART_MASK_ADDR      32'h0000_000f
`define RAM_BASE_ADDR       32'h4000_0000
`define RAM_BASE            32'h4000_0000
`define RAM_MASK_ADDR       32'h0007_ffff
`define TIMER_BASE_ADDR     32'h3000_0000
`define TIMER_MASK_ADDR     32'h0000_000f


//-------�nbellek Denetleyiciler----------
`define L1_BLOK_BIT 32    
`define L1B_SATIR   256
`define L1B_YOL     2  
`define L1V_SATIR   256
`define L1V_YOL     2
`define L1_BOYUT    (`L1_BLOK_BIT * `L1B_SATIR * `L1B_YOL) + (`L1_BLOK_BIT * `L1V_SATIR * `L1V_YOL) // Teknofest 2022-2023 icin 4KB olmali
`define L1_ONBELLEK_GECIKME 1 // Denetleyici gecikmesi degil, SRAM/BRAM gecikmesi

`define ADRES_OZEL_DAGITIM
`define ADRES_BUYRUK_OZEL_BIT 0
`define ADRES_VERI_OZEL_BIT   0
`define ADRES_BYTE_BIT      2 // Veriyi byte adreslemek icin gereken bit
`define ADRES_BYTE_OFFSET   0 // ADRES_BYTE ilk bitine erismek icin gereken kaydirma
`define ADRES_SATIR_BIT     8 // Satirlari indexlemek icin gereken bit
`define ADRES_SATIR_OFFSET  (`ADRES_BYTE_OFFSET + `ADRES_BYTE_BIT) // ADRES_SATIR ilk bitine erismek icin gereken kaydirma
`define ADRES_ETIKET_BIT    (`ADRES_BIT - `ADRES_SATIR_BIT - `ADRES_BYTE_BIT) // Adresin kalan kismi
`define ADRES_ETIKET_OFFSET (`ADRES_SATIR_OFFSET + `ADRES_SATIR_BIT) // Adresin kalan kismi

`define L1_BLOK_BYTE (`L1_BLOK_BIT / 8)

// ----Yard�mc� Tan�mlamalar----
`define ALL_ONES_256        256'hFFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF
`define ALL_ONES_128        128'hFFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF_FFFF
`define ALL_ONES_64          64'hFFFF_FFFF_FFFF_FFFF
`define ALL_ONES_32          32'hFFFF_FFFF

// ----Maskeleme ��in Yard�mc� Tan�mlar----
`define NOP_MASKE           4'b0000  // B�yle mi olmal� ?

`define BYTE_MAKSE_0        4'b0001
`define BYTE_MAKSE_1        4'b0010
`define BYTE_MAKSE_2        4'b0100
`define BYTE_MAKSE_3        4'b1000

`define HALF_WORD_MASKE_0   4'b0011
`define HALF_WORD_MASKE_1   4'b0110  // Bu eri�imi yapabildi�iniz varsayd�k
`define HALF_WORD_MASKE_2   4'b1100

`define WORD_MASKE          4'b1111